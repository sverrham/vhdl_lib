--==========================================================================================
-- This VVC was generated with UVVM VVC Generator
--==========================================================================================


context vvc_context is
  library vip_vld_rdy;
  use vip_vld_rdy.transaction_pkg.all;
  use vip_vld_rdy.vvc_methods_pkg.all;
  use vip_vld_rdy.td_vvc_framework_common_methods_pkg.all;
  use vip_vld_rdy.vld_rdy_bfm_pkg.all;
end context;
