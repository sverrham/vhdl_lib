
library ieee;
use ieee.std_logic_1164.all;

package com_pkg is

	type vec8_array is array (integer range <>) of std_logic_vector(7 downto 0);

end package com_pkg;
 